package types;

    // Common
    typedef logic[ 7:0] u8_t;
    typedef logic[31:0] u32_t;

    // Memory
    typedef logic[3:0] wrstb_t;

endpackage

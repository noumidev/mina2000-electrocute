/*
 * MINA2000 "ElectroCute" is the MINAv2 reference implementation.
 * Copyright (C) 2025  noumidev
 */

module top(
    input logic clk,
    input logic rst_n
);

endmodule
